library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.vga_controller_cfg.all;

architecture arch_vga_mode of tlv_pc_ifc is

   signal vga_mode : std_logic_vector(60 downto 0);

   signal red : std_logic_vector(2 downto 0);
   signal green : std_logic_vector(2 downto 0);
   signal blue : std_logic_vector(2 downto 0);
   signal rgb : std_logic_vector(8 downto 0);
   signal rgbf : std_logic_vector(8 downto 0);
   signal vgaRow : std_logic_vector(11 downto 0);
   signal vgaCol : std_logic_vector(11 downto 0);

   signal output : std_logic; -- prepinani vystupu stopky / hodiny

   signal enable : std_logic;
   signal timeReset : std_logic;
   signal timeSet : std_logic;

   signal key : std_logic_vector(15 downto 0);
   signal digit_clr : std_logic;
   signal digit_idx : integer range 0 to 10 := 0; -- index cislice
   signal rom_col : integer range 0 to 32; -- sloupec v ROM pameti
   signal en_1MHz, en_1Hz, en_50Hz : std_logic;

   signal sec_sclk_0, sec_sclk_1, hour_sclk_0, hour_sclk_1, min_sclk_0, min_sclk_1 : integer range 0 to 9;
   signal sec_clk_0, sec_clk_1, hour_clk_0, hour_clk_1, min_clk_0, min_clk_1 : integer range 0 to 9;

   type memory is array(0 to 16*11-1) of std_logic_vector(0 to 63);
   signal number: memory :=  ("0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              (others => '0'),
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              (others => '0'),
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111110000000000000000000000000000000000000",
                              "0000000000000000000011111110000000000000000000000000000000000000",
                              "0000000000000000000011111110000000000000000000000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              (others => '0'),
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              (others => '0'),
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              (others => '0'),
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111110000000000000000000000000000000000000",
                              "0000000000000000000011111110000000000000000000000000000000000000",
                              "0000000000000000000011111110000000000000000000000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              (others => '0'),
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111110000000000000000000000000000000000000",
                              "0000000000000000000011111110000000000000000000000000000000000000",
                              "0000000000000000000011111110000000000000000000000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              (others => '0'),
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              (others => '0'),
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              (others => '0'),
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111110000000000111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000000000000000000000111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              "0000000000000000000011111111111111111111111100000000000000000000",
                              (others => '0'),
                              "0000000000000000000000000001111111111000000000000000000000000000",
                              "0000000000000000000000000001111111111000000000000000000000000000",
                              "0000000000000000000000000001111111111000000000000000000000000000",
                              "0000000000000000000000000001111111111000000000000000000000000000",
                              "0000000000000000000000000001111111111000000000000000000000000000",
                              "0000000000000000000000000000000000000000000000000000000000000000",
                              "0000000000000000000000000000000000000000000000000000000000000000",
                              "0000000000000000000000000000000000000000000000000000000000000000",
                              "0000000000000000000000000000000000000000000000000000000000000000",
                              "0000000000000000000000000000000000000000000000000000000000000000",
                              "0000000000000000000000000001111111111000000000000000000000000000",
                              "0000000000000000000000000001111111111000000000000000000000000000",
                              "0000000000000000000000000001111111111000000000000000000000000000",
                              "0000000000000000000000000001111111111000000000000000000000000000",
                              "0000000000000000000000000001111111111000000000000000000000000000",
                              (others => '0'));

begin

  gen_1mhz: entity work.engen
     generic map (MAXVALUE => 25)
     port map (
        CLK => CLK,
        ENABLE => '1',
        EN => en_1MHz
     );

  gen_2hz: entity work.engen
     generic map (MAXVALUE => 1000000)
     port map (
        CLK => CLK,
        ENABLE => en_1MHz,
        EN => en_1Hz
     );

  time_stopclock_conversion : entity work.time_stopclock_generator
     port map (
        CLK => CLK,
        CLK_1Hz => en_1Hz,
        time_enable => enable,
        time_reset => timeReset,
        hour_sclk_0 => hour_sclk_0,
        hour_sclk_1 => hour_sclk_1,
        minute_sclk_0 => min_sclk_0,
        minute_sclk_1 => min_sclk_1,
        second_sclk_0 => sec_sclk_0,
        second_sclk_1 => sec_sclk_1
     );

  time_clock_conversion : entity work.time_clock_generator
     port map (
        CLK => CLK,
        CLK_1Hz => en_1Hz,
        time_set => timeSet,
        hour_clk_0 => hour_clk_0,
        hour_clk_1 => hour_clk_1,
        minute_clk_0 => min_clk_0,
        minute_clk_1 => min_clk_1,
        second_clk_0 => sec_clk_0,
        second_clk_1 => sec_clk_1
     );

   keyboard: entity keyboard_controller_high
      port map (
         CLK => CLK,
         KB_KIN => KIN,
         KB_KOUT => KOUT,
         DATA_OUT => KEY
      );

   fsm: entity work.fsm
      port map (
         CLK => CLK,
         KEY => KEY,
         ENABLE => enable,
         OUTPUT => output,
         RESET => timeReset
      );

   -- pripojeny VGA radic
   vga: entity work.vga_controller(arch_vga_controller)
      port map (
         CLK    => CLK,
         RST    => RESET,
         ENABLE => '1',
         MODE   => vga_mode,
         -- signaly rgb, column, row
         DATA_RED    => red,
         DATA_GREEN  => green,
         DATA_BLUE   => blue,
         ADDR_COLUMN => vgaCol,
         ADDR_ROW    => vgaRow,
         -- pripojeno na VGA rozhrani
         VGA_RED   => RED_V,
         VGA_GREEN => GREEN_V,
         VGA_BLUE  => BLUE_V,
         VGA_HSYNC => HSYNC_V,
         VGA_VSYNC => VSYNC_V
      );

   -- Set graphical mode (640x480, 60 Hz refresh)
   setmode(r640x480x60, vga_mode);

   -- nacteni cislic a separatoru
   process(CLK)
   begin
     if (output = '0') then
       -- zobrazi cas pro stopky (stopclock)
       if (vgaRow(11 downto 4) = "00010000") then
         if (vgaCol(11 downto 5) = "0001000") then
            digit_idx <= hour_sclk_0;
         elsif (vgaCol(11 downto 5) = "0001001") then
            digit_idx <= hour_sclk_1;
         elsif (vgaCol(11 downto 5) = "0001010") then
            digit_idx <= 10; -- separator
         elsif (vgaCol(11 downto 5) = "0001011") then
            digit_idx <= min_sclk_0;
         elsif (vgaCol(11 downto 5) = "0001100") then
            digit_idx <= min_sclk_1;
         elsif (vgaCol(11 downto 5) = "0001101") then
            digit_idx <= 10; -- separator
         elsif (vgaCol(11 downto 5) = "0001110") then
            digit_idx <= sec_sclk_0;
         elsif (vgaCol(11 downto 5) = "0001111") then
            digit_idx <= sec_sclk_1;
         end if;
       end if;
     else
       -- zobrazi cas pro hodiny (clock)
       if (vgaRow(11 downto 4) = "00010000") then
         if (vgaCol(11 downto 5) = "0001000") then
            digit_idx <= hour_clk_0;
         elsif (vgaCol(11 downto 5) = "0001001") then
            digit_idx <= hour_clk_1;
         elsif (vgaCol(11 downto 5) = "0001010") then
            digit_idx <= 10; -- separator
         elsif (vgaCol(11 downto 5) = "0001011") then
            digit_idx <= min_clk_0;
         elsif (vgaCol(11 downto 5) = "0001100") then
            digit_idx <= min_clk_1;
         elsif (vgaCol(11 downto 5) = "0001101") then
            digit_idx <= 10; -- separator
         elsif (vgaCol(11 downto 5) = "0001110") then
            digit_idx <= sec_clk_0;
         elsif (vgaCol(11 downto 5) = "0001111") then
            digit_idx <= sec_clk_1;
         end if;
       end if;
     end if;
   end process;

   rom_col <= conv_integer(vgaCol(4 downto 0)) * 2;
   digit_clr <= number(digit_idx*16 + conv_integer(vgaRow(4 downto 0)))(rom_col); -- posun cisla

   -- barva vystupu
   rgb <= "000" & "111" & "000" when digit_clr = '1' and output = '0' else -- stopky
          "111" & "000" & "000" when digit_clr = '1' and output = '1' else -- hodiny
          "000" & "000" & "000";


   -- funkce ze ktere se naplnuji rgb
   rgbf <= rgb when ((vgaCol(11 downto 5) = "0001000") and (vgaRow(11 downto 4) = "00010000")) or
                    ((vgaCol(11 downto 5) = "0001001") and (vgaRow(11 downto 4) = "00010000")) or
                    ((vgaCol(11 downto 5) = "0001010") and (vgaRow(11 downto 4) = "00010000")) or
                    ((vgaCol(11 downto 5) = "0001011") and (vgaRow(11 downto 4) = "00010000")) or
                    ((vgaCol(11 downto 5) = "0001100") and (vgaRow(11 downto 4) = "00010000")) or
                    ((vgaCol(11 downto 5) = "0001101") and (vgaRow(11 downto 4) = "00010000")) or
                    ((vgaCol(11 downto 5) = "0001110") and (vgaRow(11 downto 4) = "00010000")) or
                    ((vgaCol(11 downto 5) = "0001111") and (vgaRow(11 downto 4) = "00010000"))
               else "000" & "000" & "000";

   -- signaly k naplneni
   red <= rgbf(8 downto 6);
   green <= rgbf(5 downto 3);
   blue <= rgbf(2 downto 0);

end arch_vga_mode;
